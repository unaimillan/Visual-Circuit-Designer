module and_gate(output y, input a, input b);
  assign #1 y = a & b;
endmodule